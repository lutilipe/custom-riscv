library IEEE;
use IEEE.STD_LOGIC_1164.all;
use ieee.numeric_std.all;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity tb_somador is
end tb_somador;

architecture teste of tb_somador is

component somador is
	port (	
		x, y 	: in std_logic_vector(31 downto 0);
		s 		: out std_logic_vector(31 downto 0)
	);
end component;

signal A, B, S: std_logic_vector(31 downto 0);
begin
	instancia_somador: somador port map(x=>A,y=>B,s=>S);

	A <= std_logic_vector(to_unsigned(2, 32)), std_logic_vector(to_unsigned(3, 32)) after 20 ns;
	B <= std_logic_vector(to_unsigned(50, 32)), std_logic_vector(to_unsigned(4, 32)) after 10 ns;
end teste;